library IEEE;
use IEEE.std_logic_1164.all;

package testbench_pkg is
   constant FILE_NAME : string := "chk_sim_sig_advanced.txt";

   constant N_TEST_WORDS : integer := 1744; 
   type t_test_words     is array (1 to N_TEST_WORDS) 
                                  of string(1 to 15);
   constant test_words : t_test_words :=
   ( 
     "03799942080#   ",
     "13799942080#   ",
     "23799942080#   ",
     "33799942080#   ",
     "43799942080#   ",
     "53799942080#   ",
     "63799942080#   ",
     "73799942080#   ",
     "83799942080#   ",
     "93799942080#   ",
     "A3799942080#   ",
     "B3799942080#   ",
     "C3799942080#   ",
     "D3799942080#   ",
     "*3799942080#   ",
     "10799942080#   ",
     "11799942080#   ",
     "12799942080#   ",
     "13799942080#   ",
     "14799942080#   ",
     "15799942080#   ",
     "16799942080#   ",
     "17799942080#   ",
     "18799942080#   ",
     "19799942080#   ",
     "1A799942080#   ",
     "1B799942080#   ",
     "1C799942080#   ",
     "1D799942080#   ",
     "1*799942080#   ",
     "13099942080#   ",
     "13199942080#   ",
     "13299942080#   ",
     "13399942080#   ",
     "13499942080#   ",
     "13599942080#   ",
     "13699942080#   ",
     "13799942080#   ",
     "13899942080#   ",
     "13999942080#   ",
     "13A99942080#   ",
     "13B99942080#   ",
     "13C99942080#   ",
     "13D99942080#   ",
     "13*99942080#   ",
     "13709942080#   ",
     "13719942080#   ",
     "13729942080#   ",
     "13739942080#   ",
     "13749942080#   ",
     "13759942080#   ",
     "13769942080#   ",
     "13779942080#   ",
     "13789942080#   ",
     "13799942080#   ",
     "137A9942080#   ",
     "137B9942080#   ",
     "137C9942080#   ",
     "137D9942080#   ",
     "137*9942080#   ",
     "13790942080#   ",
     "13791942080#   ",
     "13792942080#   ",
     "13793942080#   ",
     "13794942080#   ",
     "13795942080#   ",
     "13796942080#   ",
     "13797942080#   ",
     "13798942080#   ",
     "13799942080#   ",
     "1379A942080#   ",
     "1379B942080#   ",
     "1379C942080#   ",
     "1379D942080#   ",
     "1379*942080#   ",
     "13799042080#   ",
     "13799142080#   ",
     "13799242080#   ",
     "13799342080#   ",
     "13799442080#   ",
     "13799542080#   ",
     "13799642080#   ",
     "13799742080#   ",
     "13799842080#   ",
     "13799942080#   ",
     "13799A42080#   ",
     "13799B42080#   ",
     "13799C42080#   ",
     "13799D42080#   ",
     "13799*42080#   ",
     "13799902080#   ",
     "13799912080#   ",
     "13799922080#   ",
     "13799932080#   ",
     "13799942080#   ",
     "13799952080#   ",
     "13799962080#   ",
     "13799972080#   ",
     "13799982080#   ",
     "13799992080#   ",
     "137999A2080#   ",
     "137999B2080#   ",
     "137999C2080#   ",
     "137999D2080#   ",
     "137999*2080#   ",
     "13799940080#   ",
     "13799941080#   ",
     "13799942080#   ",
     "13799943080#   ",
     "13799944080#   ",
     "13799945080#   ",
     "13799946080#   ",
     "13799947080#   ",
     "13799948080#   ",
     "13799949080#   ",
     "1379994A080#   ",
     "1379994B080#   ",
     "1379994C080#   ",
     "1379994D080#   ",
     "1379994*080#   ",
     "13799942080#   ",
     "13799942180#   ",
     "13799942280#   ",
     "13799942380#   ",
     "13799942480#   ",
     "13799942580#   ",
     "13799942680#   ",
     "13799942780#   ",
     "13799942880#   ",
     "13799942980#   ",
     "13799942A80#   ",
     "13799942B80#   ",
     "13799942C80#   ",
     "13799942D80#   ",
     "13799942*80#   ",
     "13799942000#   ",
     "13799942010#   ",
     "13799942020#   ",
     "13799942030#   ",
     "13799942040#   ",
     "13799942050#   ",
     "13799942060#   ",
     "13799942070#   ",
     "13799942080#   ",
     "13799942090#   ",
     "137999420A0#   ",
     "137999420B0#   ",
     "137999420C0#   ",
     "137999420D0#   ",
     "137999420*0#   ",
     "13799942080#   ",
     "13799942081#   ",
     "13799942082#   ",
     "13799942083#   ",
     "13799942084#   ",
     "13799942085#   ",
     "13799942086#   ",
     "13799942087#   ",
     "13799942088#   ",
     "13799942089#   ",
     "1379994208A#   ",
     "1379994208B#   ",
     "1379994208C#   ",
     "1379994208D#   ",
     "1379994208*#   ",
     "00#            ",
     "01#            ",
     "02#            ",
     "03#            ",
     "04#            ",
     "05#            ",
     "06#            ",
     "07#            ",
     "08#            ",
     "09#            ",
     "0A#            ",
     "0B#            ",
     "0C#            ",
     "0D#            ",
     "0*#            ",
     "0#             ",
     "10#            ",
     "11#            ",
     "12#            ",
     "13#            ",
     "14#            ",
     "15#            ",
     "16#            ",
     "17#            ",
     "18#            ",
     "19#            ",
     "1A#            ",
     "1B#            ",
     "1C#            ",
     "1D#            ",
     "1*#            ",
     "1#             ",
     "20#            ",
     "21#            ",
     "22#            ",
     "23#            ",
     "24#            ",
     "25#            ",
     "26#            ",
     "27#            ",
     "28#            ",
     "29#            ",
     "2A#            ",
     "2B#            ",
     "2C#            ",
     "2D#            ",
     "2*#            ",
     "2#             ",
     "30#            ",
     "31#            ",
     "32#            ",
     "33#            ",
     "34#            ",
     "35#            ",
     "36#            ",
     "37#            ",
     "38#            ",
     "39#            ",
     "3A#            ",
     "3B#            ",
     "3C#            ",
     "3D#            ",
     "3*#            ",
     "3#             ",
     "40#            ",
     "41#            ",
     "42#            ",
     "43#            ",
     "44#            ",
     "45#            ",
     "46#            ",
     "47#            ",
     "48#            ",
     "49#            ",
     "4A#            ",
     "4B#            ",
     "4C#            ",
     "4D#            ",
     "4*#            ",
     "4#             ",
     "50#            ",
     "51#            ",
     "52#            ",
     "53#            ",
     "54#            ",
     "55#            ",
     "56#            ",
     "57#            ",
     "58#            ",
     "59#            ",
     "5A#            ",
     "5B#            ",
     "5C#            ",
     "5D#            ",
     "5*#            ",
     "5#             ",
     "60#            ",
     "61#            ",
     "62#            ",
     "63#            ",
     "64#            ",
     "65#            ",
     "66#            ",
     "67#            ",
     "68#            ",
     "69#            ",
     "6A#            ",
     "6B#            ",
     "6C#            ",
     "6D#            ",
     "6*#            ",
     "6#             ",
     "70#            ",
     "71#            ",
     "72#            ",
     "73#            ",
     "74#            ",
     "75#            ",
     "76#            ",
     "77#            ",
     "78#            ",
     "79#            ",
     "7A#            ",
     "7B#            ",
     "7C#            ",
     "7D#            ",
     "7*#            ",
     "7#             ",
     "80#            ",
     "81#            ",
     "82#            ",
     "83#            ",
     "84#            ",
     "85#            ",
     "86#            ",
     "87#            ",
     "88#            ",
     "89#            ",
     "8A#            ",
     "8B#            ",
     "8C#            ",
     "8D#            ",
     "8*#            ",
     "8#             ",
     "90#            ",
     "91#            ",
     "92#            ",
     "93#            ",
     "94#            ",
     "95#            ",
     "96#            ",
     "97#            ",
     "98#            ",
     "99#            ",
     "9A#            ",
     "9B#            ",
     "9C#            ",
     "9D#            ",
     "9*#            ",
     "9#             ",
     "A0#            ",
     "A1#            ",
     "A2#            ",
     "A3#            ",
     "A4#            ",
     "A5#            ",
     "A6#            ",
     "A7#            ",
     "A8#            ",
     "A9#            ",
     "AA#            ",
     "AB#            ",
     "AC#            ",
     "AD#            ",
     "A*#            ",
     "A#             ",
     "B0#            ",
     "B1#            ",
     "B2#            ",
     "B3#            ",
     "B4#            ",
     "B5#            ",
     "B6#            ",
     "B7#            ",
     "B8#            ",
     "B9#            ",
     "BA#            ",
     "BB#            ",
     "BC#            ",
     "BD#            ",
     "B*#            ",
     "B#             ",
     "C0#            ",
     "C1#            ",
     "C2#            ",
     "C3#            ",
     "C4#            ",
     "C5#            ",
     "C6#            ",
     "C7#            ",
     "C8#            ",
     "C9#            ",
     "CA#            ",
     "CB#            ",
     "CC#            ",
     "CD#            ",
     "C*#            ",
     "C#             ",
     "D0#            ",
     "D1#            ",
     "D2#            ",
     "D3#            ",
     "D4#            ",
     "D5#            ",
     "D6#            ",
     "D7#            ",
     "D8#            ",
     "D9#            ",
     "DA#            ",
     "DB#            ",
     "DC#            ",
     "DD#            ",
     "D*#            ",
     "D#             ",
     "*0#            ",
     "*1#            ",
     "*2#            ",
     "*3#            ",
     "*4#            ",
     "*5#            ",
     "*6#            ",
     "*7#            ",
     "*8#            ",
     "*9#            ",
     "*A#            ",
     "*B#            ",
     "*C#            ",
     "*D#            ",
     "**#            ",
     "*#             ",
     "13799942000#   ",
     "13799942001#   ",
     "13799942002#   ",
     "13799942003#   ",
     "13799942004#   ",
     "13799942005#   ",
     "13799942006#   ",
     "13799942007#   ",
     "13799942008#   ",
     "13799942009#   ",
     "1379994200A#   ",
     "1379994200B#   ",
     "1379994200C#   ",
     "1379994200D#   ",
     "1379994200*#   ",
     "1379994200#    ",
     "13799942010#   ",
     "13799942011#   ",
     "13799942012#   ",
     "13799942013#   ",
     "13799942014#   ",
     "13799942015#   ",
     "13799942016#   ",
     "13799942017#   ",
     "13799942018#   ",
     "13799942019#   ",
     "1379994201A#   ",
     "1379994201B#   ",
     "1379994201C#   ",
     "1379994201D#   ",
     "1379994201*#   ",
     "1379994201#    ",
     "13799942020#   ",
     "13799942021#   ",
     "13799942022#   ",
     "13799942023#   ",
     "13799942024#   ",
     "13799942025#   ",
     "13799942026#   ",
     "13799942027#   ",
     "13799942028#   ",
     "13799942029#   ",
     "1379994202A#   ",
     "1379994202B#   ",
     "1379994202C#   ",
     "1379994202D#   ",
     "1379994202*#   ",
     "1379994202#    ",
     "13799942030#   ",
     "13799942031#   ",
     "13799942032#   ",
     "13799942033#   ",
     "13799942034#   ",
     "13799942035#   ",
     "13799942036#   ",
     "13799942037#   ",
     "13799942038#   ",
     "13799942039#   ",
     "1379994203A#   ",
     "1379994203B#   ",
     "1379994203C#   ",
     "1379994203D#   ",
     "1379994203*#   ",
     "1379994203#    ",
     "13799942040#   ",
     "13799942041#   ",
     "13799942042#   ",
     "13799942043#   ",
     "13799942044#   ",
     "13799942045#   ",
     "13799942046#   ",
     "13799942047#   ",
     "13799942048#   ",
     "13799942049#   ",
     "1379994204A#   ",
     "1379994204B#   ",
     "1379994204C#   ",
     "1379994204D#   ",
     "1379994204*#   ",
     "1379994204#    ",
     "13799942050#   ",
     "13799942051#   ",
     "13799942052#   ",
     "13799942053#   ",
     "13799942054#   ",
     "13799942055#   ",
     "13799942056#   ",
     "13799942057#   ",
     "13799942058#   ",
     "13799942059#   ",
     "1379994205A#   ",
     "1379994205B#   ",
     "1379994205C#   ",
     "1379994205D#   ",
     "1379994205*#   ",
     "1379994205#    ",
     "13799942060#   ",
     "13799942061#   ",
     "13799942062#   ",
     "13799942063#   ",
     "13799942064#   ",
     "13799942065#   ",
     "13799942066#   ",
     "13799942067#   ",
     "13799942068#   ",
     "13799942069#   ",
     "1379994206A#   ",
     "1379994206B#   ",
     "1379994206C#   ",
     "1379994206D#   ",
     "1379994206*#   ",
     "1379994206#    ",
     "13799942070#   ",
     "13799942071#   ",
     "13799942072#   ",
     "13799942073#   ",
     "13799942074#   ",
     "13799942075#   ",
     "13799942076#   ",
     "13799942077#   ",
     "13799942078#   ",
     "13799942079#   ",
     "1379994207A#   ",
     "1379994207B#   ",
     "1379994207C#   ",
     "1379994207D#   ",
     "1379994207*#   ",
     "1379994207#    ",
     "13799942080#   ",
     "13799942081#   ",
     "13799942082#   ",
     "13799942083#   ",
     "13799942084#   ",
     "13799942085#   ",
     "13799942086#   ",
     "13799942087#   ",
     "13799942088#   ",
     "13799942089#   ",
     "1379994208A#   ",
     "1379994208B#   ",
     "1379994208C#   ",
     "1379994208D#   ",
     "1379994208*#   ",
     "1379994208#    ",
     "13799942090#   ",
     "13799942091#   ",
     "13799942092#   ",
     "13799942093#   ",
     "13799942094#   ",
     "13799942095#   ",
     "13799942096#   ",
     "13799942097#   ",
     "13799942098#   ",
     "13799942099#   ",
     "1379994209A#   ",
     "1379994209B#   ",
     "1379994209C#   ",
     "1379994209D#   ",
     "1379994209*#   ",
     "1379994209#    ",
     "137999420A0#   ",
     "137999420A1#   ",
     "137999420A2#   ",
     "137999420A3#   ",
     "137999420A4#   ",
     "137999420A5#   ",
     "137999420A6#   ",
     "137999420A7#   ",
     "137999420A8#   ",
     "137999420A9#   ",
     "137999420AA#   ",
     "137999420AB#   ",
     "137999420AC#   ",
     "137999420AD#   ",
     "137999420A*#   ",
     "137999420A#    ",
     "137999420B0#   ",
     "137999420B1#   ",
     "137999420B2#   ",
     "137999420B3#   ",
     "137999420B4#   ",
     "137999420B5#   ",
     "137999420B6#   ",
     "137999420B7#   ",
     "137999420B8#   ",
     "137999420B9#   ",
     "137999420BA#   ",
     "137999420BB#   ",
     "137999420BC#   ",
     "137999420BD#   ",
     "137999420B*#   ",
     "137999420B#    ",
     "137999420C0#   ",
     "137999420C1#   ",
     "137999420C2#   ",
     "137999420C3#   ",
     "137999420C4#   ",
     "137999420C5#   ",
     "137999420C6#   ",
     "137999420C7#   ",
     "137999420C8#   ",
     "137999420C9#   ",
     "137999420CA#   ",
     "137999420CB#   ",
     "137999420CC#   ",
     "137999420CD#   ",
     "137999420C*#   ",
     "137999420C#    ",
     "137999420D0#   ",
     "137999420D1#   ",
     "137999420D2#   ",
     "137999420D3#   ",
     "137999420D4#   ",
     "137999420D5#   ",
     "137999420D6#   ",
     "137999420D7#   ",
     "137999420D8#   ",
     "137999420D9#   ",
     "137999420DA#   ",
     "137999420DB#   ",
     "137999420DC#   ",
     "137999420DD#   ",
     "137999420D*#   ",
     "137999420D#    ",
     "137999420*0#   ",
     "137999420*1#   ",
     "137999420*2#   ",
     "137999420*3#   ",
     "137999420*4#   ",
     "137999420*5#   ",
     "137999420*6#   ",
     "137999420*7#   ",
     "137999420*8#   ",
     "137999420*9#   ",
     "137999420*A#   ",
     "137999420*B#   ",
     "137999420*C#   ",
     "137999420*D#   ",
     "137999420**#   ",
     "137999420*#    ",
     "013799942080#  ",
     "113799942080#  ",
     "213799942080#  ",
     "313799942080#  ",
     "413799942080#  ",
     "513799942080#  ",
     "613799942080#  ",
     "713799942080#  ",
     "813799942080#  ",
     "913799942080#  ",
     "A13799942080#  ",
     "B13799942080#  ",
     "C13799942080#  ",
     "D13799942080#  ",
     "*13799942080#  ",
     "103799942080#  ",
     "113799942080#  ",
     "123799942080#  ",
     "133799942080#  ",
     "143799942080#  ",
     "153799942080#  ",
     "163799942080#  ",
     "173799942080#  ",
     "183799942080#  ",
     "193799942080#  ",
     "1A3799942080#  ",
     "1B3799942080#  ",
     "1C3799942080#  ",
     "1D3799942080#  ",
     "1*3799942080#  ",
     "130799942080#  ",
     "131799942080#  ",
     "132799942080#  ",
     "133799942080#  ",
     "134799942080#  ",
     "135799942080#  ",
     "136799942080#  ",
     "137799942080#  ",
     "138799942080#  ",
     "139799942080#  ",
     "13A799942080#  ",
     "13B799942080#  ",
     "13C799942080#  ",
     "13D799942080#  ",
     "13*799942080#  ",
     "137099942080#  ",
     "137199942080#  ",
     "137299942080#  ",
     "137399942080#  ",
     "137499942080#  ",
     "137599942080#  ",
     "137699942080#  ",
     "137799942080#  ",
     "137899942080#  ",
     "137999942080#  ",
     "137A99942080#  ",
     "137B99942080#  ",
     "137C99942080#  ",
     "137D99942080#  ",
     "137*99942080#  ",
     "137909942080#  ",
     "137919942080#  ",
     "137929942080#  ",
     "137939942080#  ",
     "137949942080#  ",
     "137959942080#  ",
     "137969942080#  ",
     "137979942080#  ",
     "137989942080#  ",
     "137999942080#  ",
     "1379A9942080#  ",
     "1379B9942080#  ",
     "1379C9942080#  ",
     "1379D9942080#  ",
     "1379*9942080#  ",
     "137990942080#  ",
     "137991942080#  ",
     "137992942080#  ",
     "137993942080#  ",
     "137994942080#  ",
     "137995942080#  ",
     "137996942080#  ",
     "137997942080#  ",
     "137998942080#  ",
     "137999942080#  ",
     "13799A942080#  ",
     "13799B942080#  ",
     "13799C942080#  ",
     "13799D942080#  ",
     "13799*942080#  ",
     "137999042080#  ",
     "137999142080#  ",
     "137999242080#  ",
     "137999342080#  ",
     "137999442080#  ",
     "137999542080#  ",
     "137999642080#  ",
     "137999742080#  ",
     "137999842080#  ",
     "137999942080#  ",
     "137999A42080#  ",
     "137999B42080#  ",
     "137999C42080#  ",
     "137999D42080#  ",
     "137999*42080#  ",
     "137999402080#  ",
     "137999412080#  ",
     "137999422080#  ",
     "137999432080#  ",
     "137999442080#  ",
     "137999452080#  ",
     "137999462080#  ",
     "137999472080#  ",
     "137999482080#  ",
     "137999492080#  ",
     "1379994A2080#  ",
     "1379994B2080#  ",
     "1379994C2080#  ",
     "1379994D2080#  ",
     "1379994*2080#  ",
     "137999420080#  ",
     "137999421080#  ",
     "137999422080#  ",
     "137999423080#  ",
     "137999424080#  ",
     "137999425080#  ",
     "137999426080#  ",
     "137999427080#  ",
     "137999428080#  ",
     "137999429080#  ",
     "13799942A080#  ",
     "13799942B080#  ",
     "13799942C080#  ",
     "13799942D080#  ",
     "13799942*080#  ",
     "137999420080#  ",
     "137999420180#  ",
     "137999420280#  ",
     "137999420380#  ",
     "137999420480#  ",
     "137999420580#  ",
     "137999420680#  ",
     "137999420780#  ",
     "137999420880#  ",
     "137999420980#  ",
     "137999420A80#  ",
     "137999420B80#  ",
     "137999420C80#  ",
     "137999420D80#  ",
     "137999420*80#  ",
     "137999420800#  ",
     "137999420810#  ",
     "137999420820#  ",
     "137999420830#  ",
     "137999420840#  ",
     "137999420850#  ",
     "137999420860#  ",
     "137999420870#  ",
     "137999420880#  ",
     "137999420890#  ",
     "1379994208A0#  ",
     "1379994208B0#  ",
     "1379994208C0#  ",
     "1379994208D0#  ",
     "1379994208*0#  ",
     "137999420800#  ",
     "137999420801#  ",
     "137999420802#  ",
     "137999420803#  ",
     "137999420804#  ",
     "137999420805#  ",
     "137999420806#  ",
     "137999420807#  ",
     "137999420808#  ",
     "137999420809#  ",
     "13799942080A#  ",
     "13799942080B#  ",
     "13799942080C#  ",
     "13799942080D#  ",
     "13799942080*#  ",
     "3799942080#    ",
     "1799942080#    ",
     "1399942080#    ",
     "1379942080#    ",
     "1379942080#    ",
     "1379942080#    ",
     "1379992080#    ",
     "1379994080#    ",
     "1379994280#    ",
     "1379994200#    ",
     "1379994208#    ",
     "#              ",
     "1#             ",
     "13#            ",
     "137#           ",
     "1379#          ",
     "13799#         ",
     "137999#        ",
     "1379994#       ",
     "13799942#      ",
     "137999420#     ",
     "1379994208#    ",
     "13799942080#   ",
     "13799942080#   ",
     "3799942080#    ",
     "799942080#     ",
     "99942080#      ",
     "9942080#       ",
     "942080#        ",
     "42080#         ",
     "2080#          ",
     "080#           ",
     "80#            ",
     "0#             ",
     "#              ",
     "03812975803#   ",
     "13812975803#   ",
     "23812975803#   ",
     "33812975803#   ",
     "43812975803#   ",
     "53812975803#   ",
     "63812975803#   ",
     "73812975803#   ",
     "83812975803#   ",
     "93812975803#   ",
     "A3812975803#   ",
     "B3812975803#   ",
     "C3812975803#   ",
     "D3812975803#   ",
     "*3812975803#   ",
     "10812975803#   ",
     "11812975803#   ",
     "12812975803#   ",
     "13812975803#   ",
     "14812975803#   ",
     "15812975803#   ",
     "16812975803#   ",
     "17812975803#   ",
     "18812975803#   ",
     "19812975803#   ",
     "1A812975803#   ",
     "1B812975803#   ",
     "1C812975803#   ",
     "1D812975803#   ",
     "1*812975803#   ",
     "13012975803#   ",
     "13112975803#   ",
     "13212975803#   ",
     "13312975803#   ",
     "13412975803#   ",
     "13512975803#   ",
     "13612975803#   ",
     "13712975803#   ",
     "13812975803#   ",
     "13912975803#   ",
     "13A12975803#   ",
     "13B12975803#   ",
     "13C12975803#   ",
     "13D12975803#   ",
     "13*12975803#   ",
     "13802975803#   ",
     "13812975803#   ",
     "13822975803#   ",
     "13832975803#   ",
     "13842975803#   ",
     "13852975803#   ",
     "13862975803#   ",
     "13872975803#   ",
     "13882975803#   ",
     "13892975803#   ",
     "138A2975803#   ",
     "138B2975803#   ",
     "138C2975803#   ",
     "138D2975803#   ",
     "138*2975803#   ",
     "13810975803#   ",
     "13811975803#   ",
     "13812975803#   ",
     "13813975803#   ",
     "13814975803#   ",
     "13815975803#   ",
     "13816975803#   ",
     "13817975803#   ",
     "13818975803#   ",
     "13819975803#   ",
     "1381A975803#   ",
     "1381B975803#   ",
     "1381C975803#   ",
     "1381D975803#   ",
     "1381*975803#   ",
     "13812075803#   ",
     "13812175803#   ",
     "13812275803#   ",
     "13812375803#   ",
     "13812475803#   ",
     "13812575803#   ",
     "13812675803#   ",
     "13812775803#   ",
     "13812875803#   ",
     "13812975803#   ",
     "13812A75803#   ",
     "13812B75803#   ",
     "13812C75803#   ",
     "13812D75803#   ",
     "13812*75803#   ",
     "13812905803#   ",
     "13812915803#   ",
     "13812925803#   ",
     "13812935803#   ",
     "13812945803#   ",
     "13812955803#   ",
     "13812965803#   ",
     "13812975803#   ",
     "13812985803#   ",
     "13812995803#   ",
     "138129A5803#   ",
     "138129B5803#   ",
     "138129C5803#   ",
     "138129D5803#   ",
     "138129*5803#   ",
     "13812970803#   ",
     "13812971803#   ",
     "13812972803#   ",
     "13812973803#   ",
     "13812974803#   ",
     "13812975803#   ",
     "13812976803#   ",
     "13812977803#   ",
     "13812978803#   ",
     "13812979803#   ",
     "1381297A803#   ",
     "1381297B803#   ",
     "1381297C803#   ",
     "1381297D803#   ",
     "1381297*803#   ",
     "13812975003#   ",
     "13812975103#   ",
     "13812975203#   ",
     "13812975303#   ",
     "13812975403#   ",
     "13812975503#   ",
     "13812975603#   ",
     "13812975703#   ",
     "13812975803#   ",
     "13812975903#   ",
     "13812975A03#   ",
     "13812975B03#   ",
     "13812975C03#   ",
     "13812975D03#   ",
     "13812975*03#   ",
     "13812975803#   ",
     "13812975813#   ",
     "13812975823#   ",
     "13812975833#   ",
     "13812975843#   ",
     "13812975853#   ",
     "13812975863#   ",
     "13812975873#   ",
     "13812975883#   ",
     "13812975893#   ",
     "138129758A3#   ",
     "138129758B3#   ",
     "138129758C3#   ",
     "138129758D3#   ",
     "138129758*3#   ",
     "13812975800#   ",
     "13812975801#   ",
     "13812975802#   ",
     "13812975803#   ",
     "13812975804#   ",
     "13812975805#   ",
     "13812975806#   ",
     "13812975807#   ",
     "13812975808#   ",
     "13812975809#   ",
     "1381297580A#   ",
     "1381297580B#   ",
     "1381297580C#   ",
     "1381297580D#   ",
     "1381297580*#   ",
     "00#            ",
     "01#            ",
     "02#            ",
     "03#            ",
     "04#            ",
     "05#            ",
     "06#            ",
     "07#            ",
     "08#            ",
     "09#            ",
     "0A#            ",
     "0B#            ",
     "0C#            ",
     "0D#            ",
     "0*#            ",
     "0#             ",
     "10#            ",
     "11#            ",
     "12#            ",
     "13#            ",
     "14#            ",
     "15#            ",
     "16#            ",
     "17#            ",
     "18#            ",
     "19#            ",
     "1A#            ",
     "1B#            ",
     "1C#            ",
     "1D#            ",
     "1*#            ",
     "1#             ",
     "20#            ",
     "21#            ",
     "22#            ",
     "23#            ",
     "24#            ",
     "25#            ",
     "26#            ",
     "27#            ",
     "28#            ",
     "29#            ",
     "2A#            ",
     "2B#            ",
     "2C#            ",
     "2D#            ",
     "2*#            ",
     "2#             ",
     "30#            ",
     "31#            ",
     "32#            ",
     "33#            ",
     "34#            ",
     "35#            ",
     "36#            ",
     "37#            ",
     "38#            ",
     "39#            ",
     "3A#            ",
     "3B#            ",
     "3C#            ",
     "3D#            ",
     "3*#            ",
     "3#             ",
     "40#            ",
     "41#            ",
     "42#            ",
     "43#            ",
     "44#            ",
     "45#            ",
     "46#            ",
     "47#            ",
     "48#            ",
     "49#            ",
     "4A#            ",
     "4B#            ",
     "4C#            ",
     "4D#            ",
     "4*#            ",
     "4#             ",
     "50#            ",
     "51#            ",
     "52#            ",
     "53#            ",
     "54#            ",
     "55#            ",
     "56#            ",
     "57#            ",
     "58#            ",
     "59#            ",
     "5A#            ",
     "5B#            ",
     "5C#            ",
     "5D#            ",
     "5*#            ",
     "5#             ",
     "60#            ",
     "61#            ",
     "62#            ",
     "63#            ",
     "64#            ",
     "65#            ",
     "66#            ",
     "67#            ",
     "68#            ",
     "69#            ",
     "6A#            ",
     "6B#            ",
     "6C#            ",
     "6D#            ",
     "6*#            ",
     "6#             ",
     "70#            ",
     "71#            ",
     "72#            ",
     "73#            ",
     "74#            ",
     "75#            ",
     "76#            ",
     "77#            ",
     "78#            ",
     "79#            ",
     "7A#            ",
     "7B#            ",
     "7C#            ",
     "7D#            ",
     "7*#            ",
     "7#             ",
     "80#            ",
     "81#            ",
     "82#            ",
     "83#            ",
     "84#            ",
     "85#            ",
     "86#            ",
     "87#            ",
     "88#            ",
     "89#            ",
     "8A#            ",
     "8B#            ",
     "8C#            ",
     "8D#            ",
     "8*#            ",
     "8#             ",
     "90#            ",
     "91#            ",
     "92#            ",
     "93#            ",
     "94#            ",
     "95#            ",
     "96#            ",
     "97#            ",
     "98#            ",
     "99#            ",
     "9A#            ",
     "9B#            ",
     "9C#            ",
     "9D#            ",
     "9*#            ",
     "9#             ",
     "A0#            ",
     "A1#            ",
     "A2#            ",
     "A3#            ",
     "A4#            ",
     "A5#            ",
     "A6#            ",
     "A7#            ",
     "A8#            ",
     "A9#            ",
     "AA#            ",
     "AB#            ",
     "AC#            ",
     "AD#            ",
     "A*#            ",
     "A#             ",
     "B0#            ",
     "B1#            ",
     "B2#            ",
     "B3#            ",
     "B4#            ",
     "B5#            ",
     "B6#            ",
     "B7#            ",
     "B8#            ",
     "B9#            ",
     "BA#            ",
     "BB#            ",
     "BC#            ",
     "BD#            ",
     "B*#            ",
     "B#             ",
     "C0#            ",
     "C1#            ",
     "C2#            ",
     "C3#            ",
     "C4#            ",
     "C5#            ",
     "C6#            ",
     "C7#            ",
     "C8#            ",
     "C9#            ",
     "CA#            ",
     "CB#            ",
     "CC#            ",
     "CD#            ",
     "C*#            ",
     "C#             ",
     "D0#            ",
     "D1#            ",
     "D2#            ",
     "D3#            ",
     "D4#            ",
     "D5#            ",
     "D6#            ",
     "D7#            ",
     "D8#            ",
     "D9#            ",
     "DA#            ",
     "DB#            ",
     "DC#            ",
     "DD#            ",
     "D*#            ",
     "D#             ",
     "*0#            ",
     "*1#            ",
     "*2#            ",
     "*3#            ",
     "*4#            ",
     "*5#            ",
     "*6#            ",
     "*7#            ",
     "*8#            ",
     "*9#            ",
     "*A#            ",
     "*B#            ",
     "*C#            ",
     "*D#            ",
     "**#            ",
     "*#             ",
     "13812975800#   ",
     "13812975801#   ",
     "13812975802#   ",
     "13812975803#   ",
     "13812975804#   ",
     "13812975805#   ",
     "13812975806#   ",
     "13812975807#   ",
     "13812975808#   ",
     "13812975809#   ",
     "1381297580A#   ",
     "1381297580B#   ",
     "1381297580C#   ",
     "1381297580D#   ",
     "1381297580*#   ",
     "1381297580#    ",
     "13812975810#   ",
     "13812975811#   ",
     "13812975812#   ",
     "13812975813#   ",
     "13812975814#   ",
     "13812975815#   ",
     "13812975816#   ",
     "13812975817#   ",
     "13812975818#   ",
     "13812975819#   ",
     "1381297581A#   ",
     "1381297581B#   ",
     "1381297581C#   ",
     "1381297581D#   ",
     "1381297581*#   ",
     "1381297581#    ",
     "13812975820#   ",
     "13812975821#   ",
     "13812975822#   ",
     "13812975823#   ",
     "13812975824#   ",
     "13812975825#   ",
     "13812975826#   ",
     "13812975827#   ",
     "13812975828#   ",
     "13812975829#   ",
     "1381297582A#   ",
     "1381297582B#   ",
     "1381297582C#   ",
     "1381297582D#   ",
     "1381297582*#   ",
     "1381297582#    ",
     "13812975830#   ",
     "13812975831#   ",
     "13812975832#   ",
     "13812975833#   ",
     "13812975834#   ",
     "13812975835#   ",
     "13812975836#   ",
     "13812975837#   ",
     "13812975838#   ",
     "13812975839#   ",
     "1381297583A#   ",
     "1381297583B#   ",
     "1381297583C#   ",
     "1381297583D#   ",
     "1381297583*#   ",
     "1381297583#    ",
     "13812975840#   ",
     "13812975841#   ",
     "13812975842#   ",
     "13812975843#   ",
     "13812975844#   ",
     "13812975845#   ",
     "13812975846#   ",
     "13812975847#   ",
     "13812975848#   ",
     "13812975849#   ",
     "1381297584A#   ",
     "1381297584B#   ",
     "1381297584C#   ",
     "1381297584D#   ",
     "1381297584*#   ",
     "1381297584#    ",
     "13812975850#   ",
     "13812975851#   ",
     "13812975852#   ",
     "13812975853#   ",
     "13812975854#   ",
     "13812975855#   ",
     "13812975856#   ",
     "13812975857#   ",
     "13812975858#   ",
     "13812975859#   ",
     "1381297585A#   ",
     "1381297585B#   ",
     "1381297585C#   ",
     "1381297585D#   ",
     "1381297585*#   ",
     "1381297585#    ",
     "13812975860#   ",
     "13812975861#   ",
     "13812975862#   ",
     "13812975863#   ",
     "13812975864#   ",
     "13812975865#   ",
     "13812975866#   ",
     "13812975867#   ",
     "13812975868#   ",
     "13812975869#   ",
     "1381297586A#   ",
     "1381297586B#   ",
     "1381297586C#   ",
     "1381297586D#   ",
     "1381297586*#   ",
     "1381297586#    ",
     "13812975870#   ",
     "13812975871#   ",
     "13812975872#   ",
     "13812975873#   ",
     "13812975874#   ",
     "13812975875#   ",
     "13812975876#   ",
     "13812975877#   ",
     "13812975878#   ",
     "13812975879#   ",
     "1381297587A#   ",
     "1381297587B#   ",
     "1381297587C#   ",
     "1381297587D#   ",
     "1381297587*#   ",
     "1381297587#    ",
     "13812975880#   ",
     "13812975881#   ",
     "13812975882#   ",
     "13812975883#   ",
     "13812975884#   ",
     "13812975885#   ",
     "13812975886#   ",
     "13812975887#   ",
     "13812975888#   ",
     "13812975889#   ",
     "1381297588A#   ",
     "1381297588B#   ",
     "1381297588C#   ",
     "1381297588D#   ",
     "1381297588*#   ",
     "1381297588#    ",
     "13812975890#   ",
     "13812975891#   ",
     "13812975892#   ",
     "13812975893#   ",
     "13812975894#   ",
     "13812975895#   ",
     "13812975896#   ",
     "13812975897#   ",
     "13812975898#   ",
     "13812975899#   ",
     "1381297589A#   ",
     "1381297589B#   ",
     "1381297589C#   ",
     "1381297589D#   ",
     "1381297589*#   ",
     "1381297589#    ",
     "138129758A0#   ",
     "138129758A1#   ",
     "138129758A2#   ",
     "138129758A3#   ",
     "138129758A4#   ",
     "138129758A5#   ",
     "138129758A6#   ",
     "138129758A7#   ",
     "138129758A8#   ",
     "138129758A9#   ",
     "138129758AA#   ",
     "138129758AB#   ",
     "138129758AC#   ",
     "138129758AD#   ",
     "138129758A*#   ",
     "138129758A#    ",
     "138129758B0#   ",
     "138129758B1#   ",
     "138129758B2#   ",
     "138129758B3#   ",
     "138129758B4#   ",
     "138129758B5#   ",
     "138129758B6#   ",
     "138129758B7#   ",
     "138129758B8#   ",
     "138129758B9#   ",
     "138129758BA#   ",
     "138129758BB#   ",
     "138129758BC#   ",
     "138129758BD#   ",
     "138129758B*#   ",
     "138129758B#    ",
     "138129758C0#   ",
     "138129758C1#   ",
     "138129758C2#   ",
     "138129758C3#   ",
     "138129758C4#   ",
     "138129758C5#   ",
     "138129758C6#   ",
     "138129758C7#   ",
     "138129758C8#   ",
     "138129758C9#   ",
     "138129758CA#   ",
     "138129758CB#   ",
     "138129758CC#   ",
     "138129758CD#   ",
     "138129758C*#   ",
     "138129758C#    ",
     "138129758D0#   ",
     "138129758D1#   ",
     "138129758D2#   ",
     "138129758D3#   ",
     "138129758D4#   ",
     "138129758D5#   ",
     "138129758D6#   ",
     "138129758D7#   ",
     "138129758D8#   ",
     "138129758D9#   ",
     "138129758DA#   ",
     "138129758DB#   ",
     "138129758DC#   ",
     "138129758DD#   ",
     "138129758D*#   ",
     "138129758D#    ",
     "138129758*0#   ",
     "138129758*1#   ",
     "138129758*2#   ",
     "138129758*3#   ",
     "138129758*4#   ",
     "138129758*5#   ",
     "138129758*6#   ",
     "138129758*7#   ",
     "138129758*8#   ",
     "138129758*9#   ",
     "138129758*A#   ",
     "138129758*B#   ",
     "138129758*C#   ",
     "138129758*D#   ",
     "138129758**#   ",
     "138129758*#    ",
     "013812975803#  ",
     "113812975803#  ",
     "213812975803#  ",
     "313812975803#  ",
     "413812975803#  ",
     "513812975803#  ",
     "613812975803#  ",
     "713812975803#  ",
     "813812975803#  ",
     "913812975803#  ",
     "A13812975803#  ",
     "B13812975803#  ",
     "C13812975803#  ",
     "D13812975803#  ",
     "*13812975803#  ",
     "103812975803#  ",
     "113812975803#  ",
     "123812975803#  ",
     "133812975803#  ",
     "143812975803#  ",
     "153812975803#  ",
     "163812975803#  ",
     "173812975803#  ",
     "183812975803#  ",
     "193812975803#  ",
     "1A3812975803#  ",
     "1B3812975803#  ",
     "1C3812975803#  ",
     "1D3812975803#  ",
     "1*3812975803#  ",
     "130812975803#  ",
     "131812975803#  ",
     "132812975803#  ",
     "133812975803#  ",
     "134812975803#  ",
     "135812975803#  ",
     "136812975803#  ",
     "137812975803#  ",
     "138812975803#  ",
     "139812975803#  ",
     "13A812975803#  ",
     "13B812975803#  ",
     "13C812975803#  ",
     "13D812975803#  ",
     "13*812975803#  ",
     "138012975803#  ",
     "138112975803#  ",
     "138212975803#  ",
     "138312975803#  ",
     "138412975803#  ",
     "138512975803#  ",
     "138612975803#  ",
     "138712975803#  ",
     "138812975803#  ",
     "138912975803#  ",
     "138A12975803#  ",
     "138B12975803#  ",
     "138C12975803#  ",
     "138D12975803#  ",
     "138*12975803#  ",
     "138102975803#  ",
     "138112975803#  ",
     "138122975803#  ",
     "138132975803#  ",
     "138142975803#  ",
     "138152975803#  ",
     "138162975803#  ",
     "138172975803#  ",
     "138182975803#  ",
     "138192975803#  ",
     "1381A2975803#  ",
     "1381B2975803#  ",
     "1381C2975803#  ",
     "1381D2975803#  ",
     "1381*2975803#  ",
     "138120975803#  ",
     "138121975803#  ",
     "138122975803#  ",
     "138123975803#  ",
     "138124975803#  ",
     "138125975803#  ",
     "138126975803#  ",
     "138127975803#  ",
     "138128975803#  ",
     "138129975803#  ",
     "13812A975803#  ",
     "13812B975803#  ",
     "13812C975803#  ",
     "13812D975803#  ",
     "13812*975803#  ",
     "138129075803#  ",
     "138129175803#  ",
     "138129275803#  ",
     "138129375803#  ",
     "138129475803#  ",
     "138129575803#  ",
     "138129675803#  ",
     "138129775803#  ",
     "138129875803#  ",
     "138129975803#  ",
     "138129A75803#  ",
     "138129B75803#  ",
     "138129C75803#  ",
     "138129D75803#  ",
     "138129*75803#  ",
     "138129705803#  ",
     "138129715803#  ",
     "138129725803#  ",
     "138129735803#  ",
     "138129745803#  ",
     "138129755803#  ",
     "138129765803#  ",
     "138129775803#  ",
     "138129785803#  ",
     "138129795803#  ",
     "1381297A5803#  ",
     "1381297B5803#  ",
     "1381297C5803#  ",
     "1381297D5803#  ",
     "1381297*5803#  ",
     "138129750803#  ",
     "138129751803#  ",
     "138129752803#  ",
     "138129753803#  ",
     "138129754803#  ",
     "138129755803#  ",
     "138129756803#  ",
     "138129757803#  ",
     "138129758803#  ",
     "138129759803#  ",
     "13812975A803#  ",
     "13812975B803#  ",
     "13812975C803#  ",
     "13812975D803#  ",
     "13812975*803#  ",
     "138129758003#  ",
     "138129758103#  ",
     "138129758203#  ",
     "138129758303#  ",
     "138129758403#  ",
     "138129758503#  ",
     "138129758603#  ",
     "138129758703#  ",
     "138129758803#  ",
     "138129758903#  ",
     "138129758A03#  ",
     "138129758B03#  ",
     "138129758C03#  ",
     "138129758D03#  ",
     "138129758*03#  ",
     "138129758003#  ",
     "138129758013#  ",
     "138129758023#  ",
     "138129758033#  ",
     "138129758043#  ",
     "138129758053#  ",
     "138129758063#  ",
     "138129758073#  ",
     "138129758083#  ",
     "138129758093#  ",
     "1381297580A3#  ",
     "1381297580B3#  ",
     "1381297580C3#  ",
     "1381297580D3#  ",
     "1381297580*3#  ",
     "138129758030#  ",
     "138129758031#  ",
     "138129758032#  ",
     "138129758033#  ",
     "138129758034#  ",
     "138129758035#  ",
     "138129758036#  ",
     "138129758037#  ",
     "138129758038#  ",
     "138129758039#  ",
     "13812975803A#  ",
     "13812975803B#  ",
     "13812975803C#  ",
     "13812975803D#  ",
     "13812975803*#  ",
     "3812975803#    ",
     "1812975803#    ",
     "1312975803#    ",
     "1382975803#    ",
     "1381975803#    ",
     "1381275803#    ",
     "1381295803#    ",
     "1381297803#    ",
     "1381297503#    ",
     "1381297583#    ",
     "1381297580#    ",
     "#              ",
     "1#             ",
     "13#            ",
     "138#           ",
     "1381#          ",
     "13812#         ",
     "138129#        ",
     "1381297#       ",
     "13812975#      ",
     "138129758#     ",
     "1381297580#    ",
     "13812975803#   ",
     "13812975803#   ",
     "3812975803#    ",
     "812975803#     ",
     "12975803#      ",
     "2975803#       ",
     "975803#        ",
     "75803#         ",
     "5803#          ",
     "803#           ",
     "03#            ",
     "3#             ",
     "#              ",
     "13799942080#   ",
     "13799942080#   ",
     "13799942080#   ",
     "13899942080#   ",
     "13819942080#   ",
     "13812942080#   ",
     "13812942080#   ",
     "13812972080#   ",
     "13812975080#   ",
     "13812975880#   ",
     "13812975800#   ",
     "13812975803#   ",
     "13812975803#   ",
     "13812975803#   ",
     "13812975803#   ",
     "13712975803#   ",
     "13792975803#   ",
     "13799975803#   ",
     "13799975803#   ",
     "13799945803#   ",
     "13799942803#   ",
     "13799942003#   ",
     "13799942083#   ",
     "13799942080#   "
   ); 

end testbench_pkg;

package body testbench_pkg is
end testbench_pkg;
