library IEEE;
use IEEE.std_logic_1164.all;

package testbench_pkg is
   constant FILE_NAME : string := "chk_sim_sig_basic.txt";

   constant N_TEST_WORDS : integer := 48; 
   type t_test_words     is array (1 to N_TEST_WORDS) 
                                  of string(1 to 15);
   constant test_words : t_test_words :=
   ( 
     "13799942080#   ",
     "1234567890*#   ",
     "13799942080#   ",
     "234567890*#    ",
     "13799942080#   ",
     "34567890*#     ",
     "13799942080#   ",
     "4567890*#      ",
     "13799942080#   ",
     "567890*#       ",
     "13799942080#   ",
     "67890*#        ",
     "13799942080#   ",
     "7890*#         ",
     "13799942080#   ",
     "890*#          ",
     "13799942080#   ",
     "90*#           ",
     "13799942080#   ",
     "0*#            ",
     "13799942080#   ",
     "*#             ",
     "13799942080#   ",
     "#              ",
     "13812975803#   ",
     "1234567890*#   ",
     "13812975803#   ",
     "234567890*#    ",
     "13812975803#   ",
     "34567890*#     ",
     "13812975803#   ",
     "4567890*#      ",
     "13812975803#   ",
     "567890*#       ",
     "13812975803#   ",
     "67890*#        ",
     "13812975803#   ",
     "7890*#         ",
     "13812975803#   ",
     "890*#          ",
     "13812975803#   ",
     "90*#           ",
     "13812975803#   ",
     "0*#            ",
     "13812975803#   ",
     "*#             ",
     "13812975803#   ",
     "#              "
   ); 

end testbench_pkg;

package body testbench_pkg is
end testbench_pkg;
